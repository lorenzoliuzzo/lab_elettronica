*** Differentiator circuit ***
.include UA741.SPI

Vin 1 0 DC 0 AC 1 
Rgen 0 1 50
C 1 2 2.27e-9
R 2 3 9.94K
XOA 0 2 10 11 3 UA741
VSP 10 0 12V
VSN 11 0 -12V

.control
ac dec 100 10 5e6

set color0 = white
set color1 = black 
set color2 = blue
plot db(v(3)) 
plot phase(v(3))
print db(v(3)) phase(v(3))
.endc

.end
